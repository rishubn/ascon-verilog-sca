//                              -*- Mode: Verilog -*-
// Filename        : config_sca.vh
// Description     : Parameters for SCA countermeasures
// Author          : Rishub Nagpal (rishub.nagpal 'at' iaik.tugraz.at, github.com/rishubn)
// Created On      : Tue Oct 31 15:26:22 2023
// Last Modified By: Rishub Nagpal 
// Last Modified On: Tue Oct 31 15:26:22 2023
// Update Count    : 0


`ifndef _config_sca_vh_
`define _config_sca_vh_
parameter unsigned SBOX_LATENCY = 1;
parameter integer NUM_SHARES = 2;
`endif
